LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY SPI IS
	GENERIC (
		SLAVE : INTEGER := 8;
		SLAVE_DATA_BITS : INTEGER := 2
	);
	PORT (
		CLK : IN STD_LOGIC;
		RESET : IN STD_LOGIC;
		MOSI : OUT STD_LOGIC;
		MISO : IN STD_LOGIC;
		CS : BUFFER STD_LOGIC_VECTOR(SLAVE - 1 DOWNTO 0);
		SCLK : BUFFER STD_LOGIC;

		BUSY : OUT STD_LOGIC;
		CLK_DIVI : IN INTEGER;
		CS_SELECT : IN INTEGER;

		EN : IN STD_LOGIC;

		CPOL : IN STD_LOGIC;
		CPHA : IN STD_LOGIC;

		DATA_WR : IN STD_LOGIC_VECTOR(SLAVE_DATA_BITS - 1 DOWNTO 0);
		DATA_RD : OUT STD_LOGIC_VECTOR(SLAVE_DATA_BITS - 1 DOWNTO 0);

		A_CON : IN STD_LOGIC

	);
END ENTITY;

ARCHITECTURE COMP OF SPI IS
	TYPE MACHINE IS (INIT, START_RD_WR);
	SIGNAL STATE : MACHINE;
	--CREAR SEÑALES PARA MANIPULARLOS
	SIGNAL S_SLAVE : INTEGER;
	SIGNAL CLK_COUNT : INTEGER; --LIMITE, DEPENDE DEL SLAVE
	SIGNAL COUNT : INTEGER;

	SIGNAL TX_DATA : STD_LOGIC_VECTOR(SLAVE_DATA_BITS - 1 DOWNTO 0);
	SIGNAL RX_DATA : STD_LOGIC_VECTOR(SLAVE_DATA_BITS - 1 DOWNTO 0);

	SIGNAL COUNT_T : INTEGER RANGE 0 TO 2 * SLAVE_DATA_BITS + 1;
	SIGNAL BIT_COUNT : INTEGER RANGE 0 TO 2 * SLAVE_DATA_BITS;

	SIGNAL BLOCK_CHANGE : STD_LOGIC;

	SIGNAL FLAG : STD_LOGIC;

BEGIN

	PROCESS (CLK, RESET)
	BEGIN
		IF (RESET = '0') THEN
			BUSY <= '0';
			DATA_RD <= (OTHERS => '0');
			CS <= (OTHERS => '1');
			STATE <= INIT;
			MOSI <= 'Z';

		ELSIF (RISING_EDGE(CLK)) THEN
			CASE STATE IS
				WHEN INIT =>
					BUSY <= '0';
					CS <= (OTHERS => '1');
					MOSI <= 'Z';
					SCLK <= CPOL;

					FLAG <= '0';

					IF (EN = '1') THEN
						BUSY <= '1';
						STATE <= START_RD_WR;
						TX_DATA <= DATA_WR;
						COUNT_T <= 0;

						BIT_COUNT <= 2 * SLAVE_DATA_BITS;
						IF (CPHA = '1') THEN
							BIT_COUNT <= 2 * SLAVE_DATA_BITS;
						ELSE
							BIT_COUNT <= 2 * SLAVE_DATA_BITS - 1;
						END IF;

						BLOCK_CHANGE <= NOT (CPHA);--INICIALIZAR LECTURA O ESCRITURA

						IF (CS_SELECT < SLAVE) THEN
							S_SLAVE <= CS_SELECT;
						ELSE
							S_SLAVE <= 0;
						END IF;

						IF (CLK_DIVI = 0) THEN
							CLK_COUNT <= 1;
							COUNT <= 1;
						ELSE
							CLK_COUNT <= CLK_DIVI;
							COUNT <= CLK_DIVI;
						END IF;

					ELSE
						STATE <= INIT;
					END IF;
				WHEN START_RD_WR =>
					BUSY <= '1';
					CS(S_SLAVE) <= '0';

					IF (COUNT = CLK_COUNT) THEN

						COUNT <= 1;
						BLOCK_CHANGE <= NOT BLOCK_CHANGE;

						IF (COUNT_T = 2 * SLAVE_DATA_BITS + 1) THEN
							COUNT_T <= 0;
						ELSE
							COUNT_T <= COUNT_T + 1;
						END IF;

						IF (COUNT_T <= 2 * SLAVE_DATA_BITS AND CS(S_SLAVE) = '0') THEN
							SCLK <= NOT SCLK;
						END IF;

						IF (COUNT_T < BIT_COUNT AND BLOCK_CHANGE = '1') THEN
							MOSI <= TX_DATA(SLAVE_DATA_BITS - 1);
							TX_DATA <= TX_DATA(SLAVE_DATA_BITS - 2 DOWNTO 0) & '0';-- peuqños error
						END IF;

						IF (COUNT_T < BIT_COUNT + 1 AND BLOCK_CHANGE = '0' AND CS(S_SLAVE) = '0') THEN
							RX_DATA <= RX_DATA(SLAVE_DATA_BITS - 2 DOWNTO 0) & MISO;
						END IF;

						IF (COUNT_T = BIT_COUNT AND A_CON = '1') THEN
							TX_DATA <= DATA_WR;
							COUNT_T <= BIT_COUNT - (2 * SLAVE_DATA_BITS - 1);
							FLAG <= '1';
						END IF;

						IF FLAG = '1' THEN
							FLAG <= '0';
							BUSY <= '0';
							DATA_RD <= RX_DATA;
						END IF;

						IF ((COUNT_T = 2 * SLAVE_DATA_BITS + 1) AND A_CON = '0') THEN
							BUSY <= '0';
							DATA_RD <= RX_DATA;
							MOSI <= 'Z';
							CS <= (OTHERS => '1');
							STATE <= INIT;
						ELSE
							STATE <= START_RD_WR;
						END IF;
					ELSE
						COUNT <= COUNT + 1;
						STATE <= START_RD_WR;
					END IF;

			END CASE;

		END IF;
	END PROCESS;
END ARCHITECTURE;