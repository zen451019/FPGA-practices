LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ADS1115 IS

END ENTITY;

ARCHITECTURE COMP OF ADS1115 IS 
BEGIN
    -- ADS1115 implementation would go here, potentially utilizing the I2C component
END ARCHITECTURE;